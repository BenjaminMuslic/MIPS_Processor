library IEEE;
use IEEE.std_logic_1164.all;


entity decoder_5t32 is

    port(i_In : in std_logic_vector(4 downto 0);
         i_En : in std_logic;
         o_Out : out std_logic_vector(31 downto 0));
end decoder_5t32;

architecture dataflow of decoder_5t32 is

begin
--when enable is 0 set output to all 0s

	o_Out <= (others => '0') when i_En = '0' else 
                 "00000000000000000000000000000000" when i_In = "00000" else
		 "00000000000000000000000000000001" when i_In = "00000" else 
		 "00000000000000000000000000000010" when i_In = "00001" else 
		 "00000000000000000000000000000100" when i_In = "00010" else 
		 "00000000000000000000000000001000" when i_In = "00011" else 
		 "00000000000000000000000000010000" when i_In = "00100" else 
		 "00000000000000000000000000100000" when i_In = "00101" else
		 "00000000000000000000000001000000" when i_In = "00110" else
		 "00000000000000000000000010000000" when i_In = "00111" else
		 "00000000000000000000000100000000" when i_In = "01000" else
		 "00000000000000000000001000000000" when i_In = "01001" else
		 "00000000000000000000010000000000" when i_In = "01010" else
		 "00000000000000000000100000000000" when i_In = "01011" else
		 "00000000000000000001000000000000" when i_In = "01100" else
		 "00000000000000000010000000000000" when i_In = "01101" else
		 "00000000000000000100000000000000" when i_In = "01110" else
		 "00000000000000001000000000000000" when i_In = "01111" else
		 "00000000000000010000000000000000" when i_In = "10000" else
		 "00000000000000100000000000000000" when i_In = "10001" else
		 "00000000000001000000000000000000" when i_In = "10010" else
		 "00000000000010000000000000000000" when i_In = "10011" else
		 "00000000000100000000000000000000" when i_In = "10100" else
		 "00000000001000000000000000000000" when i_In = "10101" else
		 "00000000010000000000000000000000" when i_In = "10110" else
		 "00000000100000000000000000000000" when i_In = "10111" else
		 "00000001000000000000000000000000" when i_In = "11000" else
		 "00000010000000000000000000000000" when i_In = "11001" else
		 "00000100000000000000000000000000" when i_In = "11010" else
		 "00001000000000000000000000000000" when i_In = "11011" else
		 "00010000000000000000000000000000" when i_In = "11100" else
		 "00100000000000000000000000000000" when i_In = "11101" else
		 "01000000000000000000000000000000" when i_In = "11110" else
		 "10000000000000000000000000000000" when i_In = "11111" else
		  (others => '0');

end dataflow;
